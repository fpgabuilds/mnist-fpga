module tb_aether_engine_example ();
  `include "../aether_constants/aether_constants.sv"
  ;

  logic clk;
  logic [23:0] cmd;
  logic [15:0] data_output;
  logic interrupt;
  logic assert_on;

  aether_engine #(
      .DataWidth(8),
      .MaxMatrixSize(28),
      .ConvEngineCount(2),
      .DenseEngineCount(4),
      .ClkRate(143_000_000)
  ) accelerator_inst (
      .clk_i(clk),
      .clk_data_i(clk),
      .instruction_i(cmd[23:20]),
      .param_1_i(cmd[19:16]),
      .param_2_i(cmd[15:0]),
      .data_o(data_output),
      .interrupt_o(interrupt),

      .sdram_clk_en_o(),
      .sdram_bank_activate_o(),
      .sdram_address_o(),
      .sdram_cs_o(),
      .sdram_row_addr_strobe_o(),
      .sdram_column_addr_strobe_o(),
      .sdram_we_o(),
      .sdram_dqm_o(),
      .sdram_dq_io(),
      .assert_on_i(assert_on),
      .dense_out_o()
  );

  // Clock generation
  integer cycle_count = 0;
  always begin
    #5 clk = ~clk;
    cycle_count = cycle_count + 1;
    if (cycle_count >= 8000) begin
      $display("Reached 4000 cycles, stopping simulation");
      $stop;
    end
  end

  // Define a task to execute a command on the positive edge of the clock
  task automatic execute_cmd(input logic [23:0] command);
    @(posedge clk);
    cmd = command;
  endtask

  initial begin
    clk = 1'b0;
    cmd = 24'b0;
    assert_on = 1'b0;

    execute_cmd({RST, RST_FULL, 16'h0000});
    execute_cmd({NOP, 4'h0, 16'h0000});
    assert_on = 1'b1;
    $display("Loading weights  : #0, time: %t", $time);
    execute_cmd({WRR, REG_MSTRT, 16'h0000});
    execute_cmd({WRR, REG_MENDD, 16'h0011});
    execute_cmd({LDW, LDW_STRT, 16'h0000});
    $display("Conv3x3 Layer: conv1  : #1, time: %t", $time);
    execute_cmd({LDW, LDW_CONT, 16'h6261});
    execute_cmd({LDW, LDW_CONT, 16'h2A63});
    execute_cmd({LDW, LDW_CONT, 16'h4023});
    execute_cmd({LDW, LDW_CONT, 16'h797A});
    execute_cmd({LDW, LDW_CONT, 16'h7078});
    execute_cmd({LDW, LDW_MOVE, 16'h0000});
    execute_cmd({LDW, LDW_CONT, 16'h7271});
    execute_cmd({LDW, LDW_CONT, 16'h232A});
    execute_cmd({LDW, LDW_CONT, 16'h6D40});
    execute_cmd({LDW, LDW_CONT, 16'h6B6C});
    execute_cmd({LDW, LDW_CONT, 16'h6577});
    execute_cmd({LDW, LDW_CONT, 16'h2A72});
    execute_cmd({LDW, LDW_CONT, 16'h4023});
    execute_cmd({LDW, LDW_CONT, 16'h6A6E});
    execute_cmd({LDW, LDW_CONT, 16'h7569});
    execute_cmd({LDW, LDW_CONT, 16'h7776});
    execute_cmd({LDW, LDW_CONT, 16'h232A});
    execute_cmd({LDW, LDW_CONT, 16'h7440});
    execute_cmd({LDW, LDW_CONT, 16'h7273});
    $display("Weight loading complete  : #2, time: %t", $time);
    execute_cmd({LIP, LIP_STRT, 16'h0000});
    execute_cmd({LIP, LIP_CONT, 16'hAAAA});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFCFF});
    execute_cmd({LIP, LIP_CONT, 16'h3CAF});
    execute_cmd({LIP, LIP_CONT, 16'hAFAA});
    execute_cmd({LIP, LIP_CONT, 16'hAFAF});
    execute_cmd({LIP, LIP_CONT, 16'hFFF1});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hF6FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFF67});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hF4FF});
    execute_cmd({LIP, LIP_CONT, 16'hC7C1});
    execute_cmd({LIP, LIP_CONT, 16'hF6FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h1204});
    execute_cmd({LIP, LIP_CONT, 16'hFFC6});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h72FF});
    execute_cmd({LIP, LIP_CONT, 16'h0E02});
    execute_cmd({LIP, LIP_CONT, 16'hFBAC});
    execute_cmd({LIP, LIP_CONT, 16'h025E});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFFC3});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hF4FF});
    execute_cmd({LIP, LIP_CONT, 16'h0772});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFF6C});
    execute_cmd({LIP, LIP_CONT, 16'h2EB6});
    execute_cmd({LIP, LIP_CONT, 16'h0203});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFF2B});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h6CFF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hDD38});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h025F});
    execute_cmd({LIP, LIP_CONT, 16'h3D71});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hB20B});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hF6FF});
    execute_cmd({LIP, LIP_CONT, 16'h0577});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hBA02});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hCBF0});
    execute_cmd({LIP, LIP_CONT, 16'hE4FA});
    execute_cmd({LIP, LIP_CONT, 16'h0236});
    execute_cmd({LIP, LIP_CONT, 16'h6302});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hAFFF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hD62E});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h02DB});
    execute_cmd({LIP, LIP_CONT, 16'h3B02});
    execute_cmd({LIP, LIP_CONT, 16'hFFDE});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hA9FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h1502});
    execute_cmd({LIP, LIP_CONT, 16'hFFD6});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h02D5});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFFB1});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h01FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h5A02});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h022C});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFFB1});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h01FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hED53});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h022C});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFFB1});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h01FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h2D02});
    execute_cmd({LIP, LIP_CONT, 16'hFFFB});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hD5FF});
    execute_cmd({LIP, LIP_CONT, 16'h091A});
    execute_cmd({LIP, LIP_CONT, 16'h0203});
    execute_cmd({LIP, LIP_CONT, 16'h6002});
    execute_cmd({LIP, LIP_CONT, 16'hFFFC});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h01FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h2E02});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h9CFF});
    execute_cmd({LIP, LIP_CONT, 16'h2D6A});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hBE0D});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h00FF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h2502});
    execute_cmd({LIP, LIP_CONT, 16'hCACA});
    execute_cmd({LIP, LIP_CONT, 16'h4BCA});
    execute_cmd({LIP, LIP_CONT, 16'h0B1B});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hFFB2});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h5CFF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h3E02});
    execute_cmd({LIP, LIP_CONT, 16'hFFE2});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hAFFF});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h1502});
    execute_cmd({LIP, LIP_CONT, 16'hE73E});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hD3FF});
    execute_cmd({LIP, LIP_CONT, 16'h022D});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hBC1A});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h1BD9});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h1407});
    execute_cmd({LIP, LIP_CONT, 16'hFFBE});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hD8FF});
    execute_cmd({LIP, LIP_CONT, 16'h022D});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'h4202});
    execute_cmd({LIP, LIP_CONT, 16'hFF8D});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'h93D4});
    execute_cmd({LIP, LIP_CONT, 16'h0202});
    execute_cmd({LIP, LIP_CONT, 16'hB14C});
    execute_cmd({LIP, LIP_CONT, 16'hE4B1});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    execute_cmd({LIP, LIP_CONT, 16'hFFFF});
    $display("Conv3x3 Layer: conv1  : #3, time: %t", $time);
    execute_cmd({WRR, REG_BCFG1, 16'h4002});
    execute_cmd({WRR, REG_BCFG2, 16'h001C});
    execute_cmd({WRR, REG_BCFG3, 16'h0400});
    $display("Conv3x3 Layer: conv1, chunk 0  : #4, time: %t", $time);
    execute_cmd({WRR, REG_MENDD, 16'h0008});
    execute_cmd({WRR, REG_MSTRT, 16'h0000});
    execute_cmd({LDW, LDW_CWGT, 16'h0000});
    execute_cmd({NOP, 4'h0, 16'h0000});
    @(posedge data_output[0]);
    $display("Waiting until memory is done  : #5, time: %t", $time);
    execute_cmd({NOP, 4'h0, 16'h0000});
    execute_cmd({WRR, REG_CPRM1, 16'h0048});
    execute_cmd({RST, RST_CONV, 16'h0000});
    execute_cmd({CNV, 4'h0, 16'h0000});
    execute_cmd({NOP, 4'h0, 16'h0000});
    $display("Waiting until convolution is done  : #6, time: %t", $time);
    @(posedge data_output[2]);
    execute_cmd({NOP, 4'h0, 16'h0000});
    $display("Conv3x3 Layer: conv1, chunk 1  : #7, time: %t", $time);
    execute_cmd({WRR, REG_MENDD, 16'h0011});
    execute_cmd({WRR, REG_MSTRT, 16'h0009});
    execute_cmd({LDW, LDW_CWGT, 16'h0000});
    execute_cmd({NOP, 4'h0, 16'h0000});
    @(posedge data_output[0]);
    $display("Waiting until memory is done  : #8, time: %t", $time);
    execute_cmd({NOP, 4'h0, 16'h0000});
    execute_cmd({WRR, REG_CPRM1, 16'h004E});
    execute_cmd({WRR, REG_MSTRT, 16'h0012});
    execute_cmd({WRR, REG_MENDD, 16'h02B5});
    execute_cmd({RST, RST_CONV, 16'h0000});
    execute_cmd({CNV, 4'h0, 16'h0000});
    execute_cmd({NOP, 4'h0, 16'h0000});
    $display("Waiting until convolution is done  : #9, time: %t", $time);
    @(posedge data_output[2]);
    execute_cmd({NOP, 4'h0, 16'h0000});
    $display("Waiting until memory is done  : #10, time: %t", $time);
    @(posedge data_output[0]);
    execute_cmd({NOP, 4'h0, 16'h0000});

    $stop;

  end
endmodule
